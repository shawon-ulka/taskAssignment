//TestBench Generation

module tb_memory;//TestBench code start

	reg  clk;
	reg [7:0] address;
	reg [7:0] write_data;
	reg  cs;
	reg  we;
	reg  oe;
	wire [7:0] read_data;
	reg  IO_pin

endmodule//TestBench code end